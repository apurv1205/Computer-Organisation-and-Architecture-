module controller_gr10(input go,input bo,input clk,output reg[2:0]f,output reg over,output reg tsw,output reg ldn,output reg tn,output reg ldm,output reg ldp,output reg ldpp,output reg tm,output reg ldout, output reg tp,output reg tpp,output reg tout,output reg tone
    );
reg [3:0] state;
initial state<=0;
always@(posedge clk)
begin
if (state==0)
   begin
	   if(go==0)
		    state<=0;
		else
          state<=1;		
	end
else if (state==1)
   begin
	   if(go==1)
		    state<=1;
		else
          state<=2;		
	end
else if (state==2)
   begin
	   if(go==0)
		    state<=2;
		else
          state<=3;		
	end
else if (state==3)
   begin
	   if(go==1)
		    state<=3;
		else
          state<=4;		
	end
else if (state==4)
   begin
	   if(go==0)
		    state<=4;
		else
          state<=5;		
	end
else if (state==5)
   begin
	   if(bo==0)
		    state<=6;
		else
          state<=10;		
	end	
else if(state==6)
   state<=7;
else if(state==7)
   state<=8;
else if(state==8)
   state<=9;
else if(state==9)
   state<=5;	
else if(state==10)
   begin
	   if(go==0)
		    state<=11;
		else
          state<=5;		
	end	
else
   state<=11;	
if(state==0)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=0;
		ldp<=0;
		ldpp<=0;
		tm<=0;
		ldout<=0;
		tp<=0;
		tpp<=0;
		tout<=0;
		tone<=0;
		f<=0;
		over<=0;
    end
if(state==1)
    begin
	   tsw<=1;
		ldn<=1;
		tn<=0;
		ldm<=0;
		ldp<=0;
		ldpp<=0;
		tm<=0;
		ldout<=0;
		tp<=0;
		tpp<=0;
		tout<=0;
		tone<=0;
		f<=2;
		over<=0;
    end	
if(state==2)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=1;
		ldm<=1;
		ldp<=0;
		ldpp<=0;
		tm<=0;
		ldout<=0;
		tp<=0;
		tpp<=0;
		tout<=0;
		tone<=1;
		f<=4;
		over<=0;
    end	
if(state==3)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=0;
		ldp<=1;
		ldpp<=0;
		tm<=0;
		ldout<=0;
		tp<=0;
		tpp<=0;
		tout<=0;
		tone<=1;
		f<=3;
		over<=0;
    end	
if(state==4)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=0;
		ldp<=0;
		ldpp<=1;
		tm<=0;
		ldout<=0;
		tp<=0;
		tpp<=0;
		tout<=0;
		tone<=1;
		f<=3;
		over<=0;
    end	
if(state==5)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=0;
		ldp<=0;
		ldpp<=0;
		tm<=1;
		ldout<=0;
		tp<=0;
		tpp<=0;
		tout<=0;
		tone<=1;
		f<=4;
		over<=0;
    end	
if(state==6)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=0;
		ldp<=0;
		ldpp<=0;
		tm<=0;
		ldout<=1;
		tp<=1;
		tpp<=1;
		tout<=0;
		tone<=0;
		f<=5;
		over<=0;
    end	
if(state==7)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=0;
		ldp<=0;
		ldpp<=1;
		tm<=0;
		ldout<=0;
		tp<=1;
		tpp<=0;
		tout<=0;
		tone<=0;
		f<=2;
		over<=0;
    end	
if(state==8)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=0;
		ldp<=1;
		ldpp<=0;
		tm<=0;
		ldout<=0;
		tp<=0;
		tpp<=0;
		tout<=1;
		tone<=0;
		f<=3;
		over<=0;
    end	
if(state==9)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=1;
		ldp<=0;
		ldpp<=0;
		tm<=1;
		ldout<=0;
		tp<=0;
		tpp<=0;
		tout<=0;
		tone<=1;
		f<=4;
		over<=0;
    end	
if(state==10)
    begin
	   tsw<=0;
		ldn<=0;
		tn<=0;
		ldm<=0;
		ldp<=0;
		ldpp<=0;
		tm<=0;
		ldout<=1;
		tp<=0;
		tpp<=0;
		tout<=0;
		tone<=0;
		f<=3;
		over<=1;
    end		 
end
endmodule
